    Mac OS X            	   2   �      �                                      ATTR���   �   �   I                  �   I  com.apple.quarantine q/0000;4b06c042;Mail;B079C538-F924-4EA5-82EF-7CA2512CE2CC|com.apple.mail 