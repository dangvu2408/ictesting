library verilog;
use verilog.vl_types.all;
entity Basic_ALU_test_top is
    generic(
        simulation_cycle: integer := 10
    );
end Basic_ALU_test_top;
